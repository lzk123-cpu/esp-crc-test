library verilog;
use verilog.vl_types.all;
entity tb_crc3 is
end tb_crc3;
